.title KiCad schematic
.include "models/NTCLE203E3103.lib"
XU1 /NTC 0 NTCLE203E3103_B0
I1 0 /NTC {ISOURCE}
.end
